library verilog;
use verilog.vl_types.all;
entity test_6r_sum is
end test_6r_sum;
