library verilog;
use verilog.vl_types.all;
entity tb_shifrator is
end tb_shifrator;
