module tb_shifrator();

reg [9:0] X;
wire [3:0] Y;

shifrator_0to9_to_bcd uut (
    .X(X),
    .Y(Y)
);

initial begin
    X = 10'b0000000001; #10;
    X = 10'b0000000010; #10;
    X = 10'b0000000100; #10;
    X = 10'b0000001000; #10;
    X = 10'b0000010000; #10;
    X = 10'b0000100000; #10;
    X = 10'b0001000000; #10;
    X = 10'b0010000000; #10;
    X = 10'b0100000000; #10;
    X = 10'b1000000000; #10;
    $stop;
end

endmodule

